architecture rtl of test_entity is
begin
  -- empty
end rtl;
