library work;
use work.core_pkg.all;

entity test_entity is
  port (clk : in std_logic);
end entity;

architecture rtl of test_entity is
begin
end architecture;
