entity simple is
end entity simple;

architecture rtl of simple is
begin
end architecture rtl;
