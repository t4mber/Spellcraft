entity test_vector is
  port (
    data_out : out std_logic_vector
  );
end entity test_vector;