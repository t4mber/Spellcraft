entity top is
  port (
    clk : in std_logic
  );
end entity top;
