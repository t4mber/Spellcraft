library ieee;
use ieee.std_logic_1164.all;

entity first_entity is
  port (clk : in std_logic);
end entity;

architecture rtl of first_entity is
begin
end architecture;

entity second_entity is
  port (rst : in std_logic);
end entity;

architecture rtl of second_entity is
begin
end architecture;
