library ieee;
use ieee.std_logic_1164.all;

entity simple_test is
  port (clk : in std_logic);
end entity;

architecture rtl of simple_test is
begin
end architecture;
