entity test_vector_params is
  port (
    data : out std_logic_vector(7 downto 0)
  );
end entity test_vector_params;
