entity test_out is
  port (
    clk : out std_logic
  );
end entity test_out;
