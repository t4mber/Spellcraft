entity test_ports is
  port (
    clk : in std_logic
  );
end entity test_ports;
