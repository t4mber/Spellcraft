library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity test_ent is
  port (
    clk : in std_logic
  );
end test_ent;

architecture rtl of test_ent is
begin
  -- empty
end architecture;
