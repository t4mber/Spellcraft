entity test_simple_out is
  port (
    q : out bit
  );
end entity test_simple_out;
