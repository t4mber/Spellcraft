entity test_vector_simple is
  port (
    data : out std_logic_vector
  );
end entity test_vector_simple;
