entity test_inout is
  port (
    data : inout bit
  );
end entity test_inout;
