library ieee;
use ieee.std_logic_1164.all;

entity test_minimal is
end test_minimal;

architecture rtl of test_minimal is
    signal s : std_logic;
begin
end architecture;
