entity my_entity is
  port (
    signal_x : out bit
  );
end entity my_entity;
