entity test_underscore is
  port (
    my_signal : out my_type
  );
end entity test_underscore;
