library ieee;
use ieee.std_logic_1164.all;

entity test_entity is
  port (
    clk : in std_logic
  );
end test_entity;

architecture rtl of test_entity is
begin
  -- empty architecture
end architecture;
